@00000000
8C 08 02 00 8C 09 02 00 00 00 00 00 01 09 40 20 
21 08 00 0B 01 09 40 22 35 08 00 10 01 09 40 26 
01 09 40 2A 01 09 40 20 11 09 FF F5 00 00 00 00 
@00000200
00 00 00 01 00 00 FF FF 
